//======================================================
// Copyright (C) 2019 By zhoucc
// All Rights Reserved
//======================================================
// Module : CTRLWEI
// Author : CC zhou
// Contact : 
// Date : 7 .1 .2019
//=======================================================
// Description : Control configuration of Weights for 48 PECs one by one;

// Ahead get GetWei(CTRLWEI_PlsFetch) and output RdyWei;

// input GetWei, produce CTRLWEI_PlsFetch activate Pipeline 1 clk;
// collect RdyWei from DISWEI, set 1 to RdyWei of NXTPEC;
//========================================================
module CTRLWEI #(
    parameter  = 
) (
    input                   clk     ,
    input                   rst_n   ,
    input 
                            ,
    output [ `NUMPEC                    - 1 : 0 ]CTRLWEIPEC_RdyWei ,//16 b
    input  [ `NUMPEC                    - 1 : 0 ]PECCTRLWEI_GetWei ,       
);
//=====================================================================================================================
// Constant Definition :
//=====================================================================================================================





//=====================================================================================================================
// Variable Definition :
//=====================================================================================================================





//=====================================================================================================================
// Logic Design :
//=====================================================================================================================

always @ ( posedge clk or negedge rst_n ) begin
    if ( ~rst_n ) begin
        DISWEIPEC_RdyWei <= ;
    end else if (  ) begin
        DISWEIPEC_RdyWei <= DISWEIPEC_RdyWei >> 1;
    end
end




//=====================================================================================================================
// Sub-Module :
//=====================================================================================================================


endmodule