//======================================================
// Copyright (C) 2019 By zhoucc
// All Rights Reserved
//======================================================
// Module : CONFIG
// Author : CC zhou
// Contact :
// Date :   8 . 1 .2019
//=======================================================
// Description :
//========================================================
`include "../include/dw_params_presim.vh"
module  CONFIG (
    input                                              clk     ,
    input                                              rst_n   ,
    output reg [ `C_LOG_2(`LENROW)           - 1 : 0 ] CFG_LenRow, // +1 is real value
    output reg [ `BLK_WIDTH                  - 1 : 0 ] CFG_DepBlk,
    output reg [ `BLK_WIDTH                  - 1 : 0 ] CFG_NumBlk,
    output reg [ `FRAME_WIDTH                - 1 : 0 ] CFG_NumFrm,
    output reg [ `PATCH_WIDTH                - 1 : 0 ] CFG_NumPat,
    output reg [ `LAYER_WIDTH                - 1 : 0 ] CFG_NumLay,
    output reg [ 5 + 1+`POOL_KERNEL_WIDTH                -1 : 0] CFG_POOL
);
//=====================================================================================================================
// Constant Definition :
//=====================================================================================================================





//=====================================================================================================================
// Variable Definition :
//=====================================================================================================================





//=====================================================================================================================
// Logic Design :
//=====================================================================================================================
always @ ( posedge clk or negedge rst_n ) begin
    if ( !rst_n ) begin
        CFG_LenRow <= 15;
        CFG_DepBlk <= 31;
        CFG_NumBlk <= 1;
        CFG_NumFrm <= 3;
        CFG_NumPat <= 0;
        CFG_NumLay <= 7;
        CFG_POOL   <={5'd8,1'd1,3'd2};
     end else begin
        CFG_LenRow <= 15;
        CFG_DepBlk <= 31;
        CFG_NumBlk <= 1;
        CFG_NumFrm <= 3;
        CFG_NumPat <= 0;
        CFG_NumLay <= 7;
        CFG_POOL   <={5'd8,1'd1,3'd2};
    end
end





//=====================================================================================================================
// Sub-Module :
//=====================================================================================================================


endmodule
